entity ULA_Logic_Unity is
  port (
    X, Y, DIN1, DIN2, DIN3: in bit;
    S0, S1, S2 in bit
  ) ;
end ULA_Logic_Unity;

architecture arch of ULA_Logic_Unity is
begin
    S0 <= 
end arch ; -- arch